module hello;
initial begin
    $display("why,yes");
end
endmodule
