library ieee;
use ieee.std_logic_1164.all;
entity hello is
end hello;
architecture sim of hello is
begin
    process
    begin
        report "i do not understand that";
        wait;
    end process;
end sim;
